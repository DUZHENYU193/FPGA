library verilog;
use verilog.vl_types.all;
entity DDS_tb is
end DDS_tb;
